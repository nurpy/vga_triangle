




module top()




endmodule

