

module top();








endmodule

